library IEEE;
use IEEE.STD_LOGIC_1164.all;
 use work.typedefs.all;
package image_files is



constant image_cloud : flappyimage :=
((0,0,0,0,0,0,127,127,0,0,0,0),
(0,0,0,0,0,0,127,127,127,0,0,0),
(0,0,0,0,0,127,127,127,127,127,0,0),
(0,0,0,0,127,127,127,127,127,127,127,0),
(0,0,0,0,127,127,127,127,127,95,127,0),
(0,0,0,127,127,127,127,127,127,95,127,127),
(0,127,127,127,127,127,127,127,127,63,127,127),
(0,127,127,127,127,127,127,127,127,63,95,127),
(127,127,127,127,127,127,127,127,127,31,127,127),
(127,127,127,127,127,127,127,127,127,63,127,127),
(127,127,127,95,127,127,127,127,127,63,127,127),
(0,0,127,127,127,127,127,127,127,63,95,127),
(0,0,127,127,127,127,127,127,127,95,127,127),
(0,0,0,0,127,127,127,127,127,127,127,127),
(0,0,0,0,127,127,127,127,127,127,127,127),
(0,0,0,0,127,127,127,127,127,127,127,0),
(0,0,0,0,0,127,127,127,127,127,127,0)
);
constant image_flappy : flappyimage :=
((0,0,0,0,0,0,35,35,0,0,0,0),
(0,0,0,0,35,35,127,125,35,0,0,0),
(0,0,0,35,63,35,127,127,35,35,0,0),
(0,0,35,63,63,35,127,127,35,55,35,0),
(0,35,63,63,63,35,127,127,35,55,35,0),
(0,35,63,63,63,35,127,125,35,55,55,35),
(35,63,63,63,63,63,35,35,55,55,55,35),
(35,63,63,63,63,63,63,63,55,55,55,35),
(35,63,35,35,35,63,63,63,35,55,55,35),
(35,35,127,127,127,35,63,35,105,35,55,35),
(35,127,127,127,127,127,35,105,35,105,35,0),
(35,127,127,127,127,127,35,105,35,105,35,0),
(0,35,127,35,35,127,35,105,35,105,35,0),
(0,0,35,127,127,127,35,105,35,105,35,0),
(0,0,0,35,35,35,35,105,35,105,35,0),
(0,0,0,0,0,0,35,105,35,35,0,0),
(0,0,0,0,0,0,0,35,0,0,0,0)
);
constant image_mount :  mountimage :=
((0,0,17,59,59,59,59,59,59,59),
(0,0,17,59,59,59,59,59,59,59),
(0,17,17,59,59,59,59,59,59,59),
(0,17,59,17,59,59,59,59,59,59),
(17,59,59,17,59,59,59,59,59,59),
(17,59,59,59,17,59,59,59,59,59),
(17,59,59,59,17,59,59,59,17,59),
(17,59,59,59,59,17,17,17,59,59),
(0,17,59,59,59,59,59,17,59,59),
(0,17,59,59,59,59,17,59,59,59),
(0,0,17,59,59,59,17,59,59,59),
(0,0,17,59,59,17,59,59,59,59),
(0,17,59,17,17,17,59,59,59,59),
(0,17,59,59,59,17,59,59,59,59),
(17,59,59,59,17,17,59,59,59,59),
(17,59,59,59,17,59,17,59,59,59),
(17,59,59,17,59,59,17,59,59,59),
(17,59,59,17,59,59,59,17,59,59),
(0,17,59,17,59,59,59,17,17,59),
(0,17,59,17,59,17,17,59,59,59),
(0,0,17,59,17,59,59,59,59,59),
(0,0,17,59,17,59,59,59,59,59),
(0,0,0,17,59,59,59,59,59,59),
(0,0,0,17,59,59,59,59,59,59),
(0,0,17,59,59,59,59,59,59,59),
(0,0,17,59,59,59,59,59,59,59)
);
constant image_build :  buildimage :=
((0,0,0,0,0,0,0,53,53,53,53,53,53,53,53,53,53,53,53,53,53),
(0,0,0,0,0,0,0,53,95,43,43,95,43,43,95,43,43,95,43,43,95),
(0,0,0,0,0,0,0,53,95,95,95,95,95,95,95,95,95,95,95,95,95),
(0,0,0,0,43,43,43,53,95,43,43,95,43,43,95,43,43,95,43,43,95),
(0,0,0,0,43,85,85,53,95,95,95,95,95,95,95,95,95,95,95,95,95),
(0,0,0,0,43,85,43,53,95,43,43,95,43,43,95,43,43,95,43,43,95),
(0,0,0,0,43,85,85,53,95,95,95,43,43,43,43,43,43,43,43,43,43),
(0,0,0,0,43,85,85,43,43,43,43,43,85,85,85,85,85,85,85,85,85),
(0,0,0,0,43,43,43,43,43,43,43,43,85,43,43,85,85,43,43,85,85),
(0,0,0,0,43,43,43,43,43,43,43,43,85,85,85,85,85,85,85,85,85),
(0,0,0,0,0,0,0,0,0,0,0,43,43,43,43,43,43,43,43,43,43),
(0,0,43,43,43,43,43,43,43,43,43,43,43,43,43,43,43,43,43,43,43),
(43,85,43,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85),
(43,85,43,85,43,43,85,43,43,85,85,43,43,85,85,43,43,85,85,43,43),
(43,85,43,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85),
(43,43,43,85,43,43,85,43,43,85,85,43,43,85,85,43,43,85,85,43,43),
(43,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85),
(43,85,43,85,43,43,85,43,43,85,85,43,43,85,85,43,43,85,85,43,43),
(43,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85,85),
(43,43,43,43,43,43,43,43,43,43,43,43,43,43,43,43,43,43,43,43,43)
);
constant image_pipe :  pipeimage :=
((35),
(83),
(83),
(91),
(91),
(123),
(125),
(125),
(125),
(125),
(125),
(123),
(91),
(91),
(83),
(83),
(51),
(49),
(49),
(41),
(41),
(41),
(41),
(35)
);
constant image_sayi :  sayiimage :=
((0,1,0,0,0,0),
(1,1,1,1,1,1),
(85,85,85,85,85,85),
(0,0,0,0,0,0),
(0,85,0,0,85,85),
(43,43,0,43,43,1),
(1,85,0,1,85,1),
(43,43,43,43,0,1),
(85,43,43,85,0,43),
(0,43,85,0,43,85),
(85,43,0,0,43,85),
(1,85,85,0,85,1),
(1,85,43,85,85,1),
(85,43,85,43,43,85),
(0,85,0,43,43,0),
(0,85,85,1,1,0),
(85,1,1,85,1,85),
(1,1,1,1,1,1),
(85,85,85,85,1,85),
(0,0,0,0,85,0),
(0,0,0,0,0,0),
(1,1,1,0,0,1),
(1,85,1,0,0,1),
(1,0,85,1,1,85),
(85,0,0,85,85,0),
(85,1,1,1,1,0),
(1,85,1,85,85,1),
(1,0,1,0,0,1),
(85,0,85,1,1,85),
(0,0,0,85,85,0),
(43,0,0,0,0,0),
(1,0,43,43,43,43),
(1,43,43,43,43,43),
(43,43,85,85,85,85),
(85,85,0,0,0,0),
(85,85,85,85,85,85),
(43,43,43,43,43,43),
(1,85,1,85,85,1),
(43,43,43,43,43,43),
(0,43,0,43,43,0),
(85,85,85,0,85,85),
(43,43,43,0,43,43),
(1,85,1,85,85,1),
(43,85,1,85,85,43),
(0,43,43,43,43,0),
(0,0,0,0,0,0),
(0,1,1,1,1,0),
(1,85,85,85,85,1),
(1,0,0,0,0,1),
(85,1,1,1,1,85)
);
constant sinlookup :  lookuptable :=(0,1144,2287,3430,4572,5712,6850,7987,9121,10252,11380,12505,13626,14742,15855,16962,18064,19161,20252,21336,22415,23486,24550,25607,26656,27697,28729,29753,30767,31772,32768,33754,34729,35693,36647,37590,38521,39441,40348,41243,42126,42995,43852,44695,45525,46341,47143,47930,48703,49461,50203,50931,51643,52339,53020,53684,54332,54963,55578,56175,56756,57319,57865,58393,58903,59396,59870,60326,60764,61183,61584,61966,62328,62672,62997,63303,63589,63856,64104,64332,64540,64729,64898,65048,65177,65287,65376,65446,65496,65526,65536,65526,65496,65446,65376,65287,65177,65048,64898,64729,64540,64332,64104,63856,63589,63303,62997,62672,62328,61966,61584,61183,60764,60326,59870,59396,58903,58393,57865,57319,56756,56175,55578,54963,54332,53684,53020,52339,51643,50931,50203,49461,48703,47930,47143,46341,45525,44695,43852,42995,42126,41243,40348,39441,38521,37590,36647,35693,34729,33754,32768,31772,30767,29753,28729,27697,26656,25607,24550,23486,22415,21336,20252,19161,18064,16962,15855,14742,13626,12505,11380,10252,9121,7987,6850,5712,4572,3430,2287,1144,0,-1144,-2287,-3430,-4572,-5712,-6850,-7987,-9121,-10252,-11380,-12505,-13626,-14742,-15855,-16962,-18064,-19161,-20252,-21336,-22415,-23486,-24550,-25607,-26656,-27697,-28729,-29753,-30767,-31772,-32768,-33754,-34729,-35693,-36647,-37590,-38521,-39441,-40348,-41243,-42126,-42995,-43852,-44695,-45525,-46341,-47143,-47930,-48703,-49461,-50203,-50931,-51643,-52339,-53020,-53684,-54332,-54963,-55578,-56175,-56756,-57319,-57865,-58393,-58903,-59396,-59870,-60326,-60764,-61183,-61584,-61966,-62328,-62672,-62997,-63303,-63589,-63856,-64104,-64332,-64540,-64729,-64898,-65048,-65177,-65287,-65376,-65446,-65496,-65526,-65536,-65526,-65496,-65446,-65376,-65287,-65177,-65048,-64898,-64729,-64540,-64332,-64104,-63856,-63589,-63303,-62997,-62672,-62328,-61966,-61584,-61183,-60764,-60326,-59870,-59396,-58903,-58393,-57865,-57319,-56756,-56175,-55578,-54963,-54332,-53684,-53020,-52339,-51643,-50931,-50203,-49461,-48703,-47930,-47143,-46341,-45525,-44695,-43852,-42995,-42126,-41243,-40348,-39441,-38521,-37590,-36647,-35693,-34729,-33754,-32768,-31772,-30767,-29753,-28729,-27697,-26656,-25607,-24550,-23486,-22415,-21336,-20252,-19161,-18064,-16962,-15855,-14742,-13626,-12505,-11380,-10252,-9121,-7987,-6850,-5712,-4572,-3430,-2287,-1144);
constant coslookup :  lookuptable :=(65536,65526,65496,65446,65376,65287,65177,65048,64898,64729,64540,64332,64104,63856,63589,63303,62997,62672,62328,61966,61584,61183,60764,60326,59870,59396,58903,58393,57865,57319,56756,56175,55578,54963,54332,53684,53020,52339,51643,50931,50203,49461,48703,47930,47143,46341,45525,44695,43852,42995,42126,41243,40348,39441,38521,37590,36647,35693,34729,33754,32768,31772,30767,29753,28729,27697,26656,25607,24550,23486,22415,21336,20252,19161,18064,16962,15855,14742,13626,12505,11380,10252,9121,7987,6850,5712,4572,3430,2287,1144,0,-1144,-2287,-3430,-4572,-5712,-6850,-7987,-9121,-10252,-11380,-12505,-13626,-14742,-15855,-16962,-18064,-19161,-20252,-21336,-22415,-23486,-24550,-25607,-26656,-27697,-28729,-29753,-30767,-31772,-32768,-33754,-34729,-35693,-36647,-37590,-38521,-39441,-40348,-41243,-42126,-42995,-43852,-44695,-45525,-46341,-47143,-47930,-48703,-49461,-50203,-50931,-51643,-52339,-53020,-53684,-54332,-54963,-55578,-56175,-56756,-57319,-57865,-58393,-58903,-59396,-59870,-60326,-60764,-61183,-61584,-61966,-62328,-62672,-62997,-63303,-63589,-63856,-64104,-64332,-64540,-64729,-64898,-65048,-65177,-65287,-65376,-65446,-65496,-65526,-65536,-65526,-65496,-65446,-65376,-65287,-65177,-65048,-64898,-64729,-64540,-64332,-64104,-63856,-63589,-63303,-62997,-62672,-62328,-61966,-61584,-61183,-60764,-60326,-59870,-59396,-58903,-58393,-57865,-57319,-56756,-56175,-55578,-54963,-54332,-53684,-53020,-52339,-51643,-50931,-50203,-49461,-48703,-47930,-47143,-46341,-45525,-44695,-43852,-42995,-42126,-41243,-40348,-39441,-38521,-37590,-36647,-35693,-34729,-33754,-32768,-31772,-30767,-29753,-28729,-27697,-26656,-25607,-24550,-23486,-22415,-21336,-20252,-19161,-18064,-16962,-15855,-14742,-13626,-12505,-11380,-10252,-9121,-7987,-6850,-5712,-4572,-3430,-2287,-1144,0,1144,2287,3430,4572,5712,6850,7987,9121,10252,11380,12505,13626,14742,15855,16962,18064,19161,20252,21336,22415,23486,24550,25607,26656,27697,28729,29753,30767,31772,32768,33754,34729,35693,36647,37590,38521,39441,40348,41243,42126,42995,43852,44695,45525,46341,47143,47930,48703,49461,50203,50931,51643,52339,53020,53684,54332,54963,55578,56175,56756,57319,57865,58393,58903,59396,59870,60326,60764,61183,61584,61966,62328,62672,62997,63303,63589,63856,64104,64332,64540,64729,64898,65048,65177,65287,65376,65446,65496,65526);
constant image_ground :  groundimage :=((41,125,59,59,17,49,83),
(41,125,59,17,17,49,83),
(41,125,17,17,17,49,83),
(41,125,17,17,17,49,83),
(41,125,17,17,59,49,83),
(41,125,17,59,59,49,83),
(41,125,59,59,59,49,83)
);
end image_files;